module invertor
 
(
input a,
output inv_a
);

assign inv_a = ~a;

endmodule